module lut_input (in,
                  out);
    input in;
    output out;
    
    assign out = in;
endmodule
