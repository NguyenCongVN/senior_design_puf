module lut_output (in,
                   out);
    input in;
    output out;
    
    assign out = in;
endmodule
